-- entidade vazia para o testbench
entity four_bits_ripple_carry_tb is
end;

architecture structural of four_bits_ripple_carry_tb is
    signal a, b, sum : bit_vector(3 downto 0);
    signal cout : bit;

begin
    entidade : entity work.four_bits_ripple_carry(structural)
    port map (a, b, sum, cout);

    estimulo_checagem : process is

        type linha_tv is record
            a, b, sum : bit_vector(3 downto 0);
            cout : bit;
        end record;

        type vetor_linha_tv is array (natural range <>) of linha_tv;

        constant tabela_verdade : vetor_linha_tv :=
        ( --  a       b       sum     cout 
            ("0000", "0000", "0000", '0'),  -- 00 + 00 = 00, overflow 0 
            ("0000", "0001", "0001", '0'),  -- 00 + 01 = 01, overflow 0 
            ("0000", "0010", "0010", '0'),  -- 00 + 02 = 02, overflow 0 
            ("0000", "0011", "0011", '0'),  -- 00 + 03 = 03, overflow 0 
            ("0000", "0100", "0100", '0'),  -- 00 + 04 = 04, overflow 0 
            ("0000", "0101", "0101", '0'),  -- 00 + 05 = 05, overflow 0 
            ("0000", "0110", "0110", '0'),  -- 00 + 06 = 06, overflow 0 
            ("0000", "0111", "0111", '0'),  -- 00 + 07 = 07, overflow 0 
            ("0000", "1000", "1000", '0'),  -- 00 + 08 = 08, overflow 0 
            ("0000", "1001", "1001", '0'),  -- 00 + 09 = 09, overflow 0 
            ("0000", "1010", "1010", '0'),  -- 00 + 10 = 10, overflow 0 
            ("0000", "1011", "1011", '0'),  -- 00 + 11 = 11, overflow 0 
            ("0000", "1100", "1100", '0'),  -- 00 + 12 = 12, overflow 0 
            ("0000", "1101", "1101", '0'),  -- 00 + 13 = 13, overflow 0 
            ("0000", "1110", "1110", '0'),  -- 00 + 14 = 14, overflow 0 
            ("0000", "1111", "1111", '0'),  -- 00 + 15 = 15, overflow 0 
            ("0001", "0000", "0001", '0'),  -- 01 + 00 = 01, overflow 0 
            ("0001", "0001", "0010", '0'),  -- 01 + 01 = 02, overflow 0 
            ("0001", "0010", "0011", '0'),  -- 01 + 02 = 03, overflow 0 
            ("0001", "0011", "0100", '0'),  -- 01 + 03 = 04, overflow 0 
            ("0001", "0100", "0101", '0'),  -- 01 + 04 = 05, overflow 0 
            ("0001", "0101", "0110", '0'),  -- 01 + 05 = 06, overflow 0 
            ("0001", "0110", "0111", '0'),  -- 01 + 06 = 07, overflow 0 
            ("0001", "0111", "1000", '0'),  -- 01 + 07 = 08, overflow 0 
            ("0001", "1000", "1001", '0'),  -- 01 + 08 = 09, overflow 0 
            ("0001", "1001", "1010", '0'),  -- 01 + 09 = 10, overflow 0 
            ("0001", "1010", "1011", '0'),  -- 01 + 10 = 11, overflow 0 
            ("0001", "1011", "1100", '0'),  -- 01 + 11 = 12, overflow 0 
            ("0001", "1100", "1101", '0'),  -- 01 + 12 = 13, overflow 0 
            ("0001", "1101", "1110", '0'),  -- 01 + 13 = 14, overflow 0 
            ("0001", "1110", "1111", '0'),  -- 01 + 14 = 15, overflow 0 
            ("0001", "1111", "0000", '1'),  -- 01 + 15 = 16, overflow 1 
            ("0010", "0000", "0010", '0'),  -- 02 + 00 = 02, overflow 0 
            ("0010", "0001", "0011", '0'),  -- 02 + 01 = 03, overflow 0 
            ("0010", "0010", "0100", '0'),  -- 02 + 02 = 04, overflow 0 
            ("0010", "0011", "0101", '0'),  -- 02 + 03 = 05, overflow 0 
            ("0010", "0100", "0110", '0'),  -- 02 + 04 = 06, overflow 0 
            ("0010", "0101", "0111", '0'),  -- 02 + 05 = 07, overflow 0 
            ("0010", "0110", "1000", '0'),  -- 02 + 06 = 08, overflow 0 
            ("0010", "0111", "1001", '0'),  -- 02 + 07 = 09, overflow 0 
            ("0010", "1000", "1010", '0'),  -- 02 + 08 = 10, overflow 0 
            ("0010", "1001", "1011", '0'),  -- 02 + 09 = 11, overflow 0 
            ("0010", "1010", "1100", '0'),  -- 02 + 10 = 12, overflow 0 
            ("0010", "1011", "1101", '0'),  -- 02 + 11 = 13, overflow 0 
            ("0010", "1100", "1110", '0'),  -- 02 + 12 = 14, overflow 0 
            ("0010", "1101", "1111", '0'),  -- 02 + 13 = 15, overflow 0 
            ("0010", "1110", "0000", '1'),  -- 02 + 14 = 16, overflow 1 
            ("0010", "1111", "0001", '1'),  -- 02 + 15 = 17, overflow 1 
            ("0011", "0000", "0011", '0'),  -- 03 + 00 = 03, overflow 0 
            ("0011", "0001", "0100", '0'),  -- 03 + 01 = 04, overflow 0 
            ("0011", "0010", "0101", '0'),  -- 03 + 02 = 05, overflow 0 
            ("0011", "0011", "0110", '0'),  -- 03 + 03 = 06, overflow 0 
            ("0011", "0100", "0111", '0'),  -- 03 + 04 = 07, overflow 0 
            ("0011", "0101", "1000", '0'),  -- 03 + 05 = 08, overflow 0 
            ("0011", "0110", "1001", '0'),  -- 03 + 06 = 09, overflow 0 
            ("0011", "0111", "1010", '0'),  -- 03 + 07 = 10, overflow 0 
            ("0011", "1000", "1011", '0'),  -- 03 + 08 = 11, overflow 0 
            ("0011", "1001", "1100", '0'),  -- 03 + 09 = 12, overflow 0 
            ("0011", "1010", "1101", '0'),  -- 03 + 10 = 13, overflow 0 
            ("0011", "1011", "1110", '0'),  -- 03 + 11 = 14, overflow 0 
            ("0011", "1100", "1111", '0'),  -- 03 + 12 = 15, overflow 0 
            ("0011", "1101", "0000", '1'),  -- 03 + 13 = 16, overflow 1 
            ("0011", "1110", "0001", '1'),  -- 03 + 14 = 17, overflow 1 
            ("0011", "1111", "0010", '1'),  -- 03 + 15 = 18, overflow 1 
            ("0100", "0000", "0100", '0'),  -- 04 + 00 = 04, overflow 0 
            ("0100", "0001", "0101", '0'),  -- 04 + 01 = 05, overflow 0 
            ("0100", "0010", "0110", '0'),  -- 04 + 02 = 06, overflow 0 
            ("0100", "0011", "0111", '0'),  -- 04 + 03 = 07, overflow 0 
            ("0100", "0100", "1000", '0'),  -- 04 + 04 = 08, overflow 0 
            ("0100", "0101", "1001", '0'),  -- 04 + 05 = 09, overflow 0 
            ("0100", "0110", "1010", '0'),  -- 04 + 06 = 10, overflow 0 
            ("0100", "0111", "1011", '0'),  -- 04 + 07 = 11, overflow 0 
            ("0100", "1000", "1100", '0'),  -- 04 + 08 = 12, overflow 0 
            ("0100", "1001", "1101", '0'),  -- 04 + 09 = 13, overflow 0 
            ("0100", "1010", "1110", '0'),  -- 04 + 10 = 14, overflow 0 
            ("0100", "1011", "1111", '0'),  -- 04 + 11 = 15, overflow 0 
            ("0100", "1100", "0000", '1'),  -- 04 + 12 = 16, overflow 1 
            ("0100", "1101", "0001", '1'),  -- 04 + 13 = 17, overflow 1 
            ("0100", "1110", "0010", '1'),  -- 04 + 14 = 18, overflow 1 
            ("0100", "1111", "0011", '1'),  -- 04 + 15 = 19, overflow 1 
            ("0101", "0000", "0101", '0'),  -- 05 + 00 = 05, overflow 0 
            ("0101", "0001", "0110", '0'),  -- 05 + 01 = 06, overflow 0 
            ("0101", "0010", "0111", '0'),  -- 05 + 02 = 07, overflow 0 
            ("0101", "0011", "1000", '0'),  -- 05 + 03 = 08, overflow 0 
            ("0101", "0100", "1001", '0'),  -- 05 + 04 = 09, overflow 0 
            ("0101", "0101", "1010", '0'),  -- 05 + 05 = 10, overflow 0 
            ("0101", "0110", "1011", '0'),  -- 05 + 06 = 11, overflow 0 
            ("0101", "0111", "1100", '0'),  -- 05 + 07 = 12, overflow 0 
            ("0101", "1000", "1101", '0'),  -- 05 + 08 = 13, overflow 0 
            ("0101", "1001", "1110", '0'),  -- 05 + 09 = 14, overflow 0 
            ("0101", "1010", "1111", '0'),  -- 05 + 10 = 15, overflow 0 
            ("0101", "1011", "0000", '1'),  -- 05 + 11 = 16, overflow 1 
            ("0101", "1100", "0001", '1'),  -- 05 + 12 = 17, overflow 1 
            ("0101", "1101", "0010", '1'),  -- 05 + 13 = 18, overflow 1 
            ("0101", "1110", "0011", '1'),  -- 05 + 14 = 19, overflow 1 
            ("0101", "1111", "0100", '1'),  -- 05 + 15 = 20, overflow 1 
            ("0110", "0000", "0110", '0'),  -- 06 + 00 = 06, overflow 0 
            ("0110", "0001", "0111", '0'),  -- 06 + 01 = 07, overflow 0 
            ("0110", "0010", "1000", '0'),  -- 06 + 02 = 08, overflow 0 
            ("0110", "0011", "1001", '0'),  -- 06 + 03 = 09, overflow 0 
            ("0110", "0100", "1010", '0'),  -- 06 + 04 = 10, overflow 0 
            ("0110", "0101", "1011", '0'),  -- 06 + 05 = 11, overflow 0 
            ("0110", "0110", "1100", '0'),  -- 06 + 06 = 12, overflow 0 
            ("0110", "0111", "1101", '0'),  -- 06 + 07 = 13, overflow 0 
            ("0110", "1000", "1110", '0'),  -- 06 + 08 = 14, overflow 0 
            ("0110", "1001", "1111", '0'),  -- 06 + 09 = 15, overflow 0 
            ("0110", "1010", "0000", '1'),  -- 06 + 10 = 16, overflow 1 
            ("0110", "1011", "0001", '1'),  -- 06 + 11 = 17, overflow 1 
            ("0110", "1100", "0010", '1'),  -- 06 + 12 = 18, overflow 1 
            ("0110", "1101", "0011", '1'),  -- 06 + 13 = 19, overflow 1 
            ("0110", "1110", "0100", '1'),  -- 06 + 14 = 20, overflow 1 
            ("0110", "1111", "0101", '1'),  -- 06 + 15 = 21, overflow 1 
            ("0111", "0000", "0111", '0'),  -- 07 + 00 = 07, overflow 0 
            ("0111", "0001", "1000", '0'),  -- 07 + 01 = 08, overflow 0 
            ("0111", "0010", "1001", '0'),  -- 07 + 02 = 09, overflow 0 
            ("0111", "0011", "1010", '0'),  -- 07 + 03 = 10, overflow 0 
            ("0111", "0100", "1011", '0'),  -- 07 + 04 = 11, overflow 0 
            ("0111", "0101", "1100", '0'),  -- 07 + 05 = 12, overflow 0 
            ("0111", "0110", "1101", '0'),  -- 07 + 06 = 13, overflow 0 
            ("0111", "0111", "1110", '0'),  -- 07 + 07 = 14, overflow 0 
            ("0111", "1000", "1111", '0'),  -- 07 + 08 = 15, overflow 0 
            ("0111", "1001", "0000", '1'),  -- 07 + 09 = 16, overflow 1 
            ("0111", "1010", "0001", '1'),  -- 07 + 10 = 17, overflow 1 
            ("0111", "1011", "0010", '1'),  -- 07 + 11 = 18, overflow 1 
            ("0111", "1100", "0011", '1'),  -- 07 + 12 = 19, overflow 1 
            ("0111", "1101", "0100", '1'),  -- 07 + 13 = 20, overflow 1 
            ("0111", "1110", "0101", '1'),  -- 07 + 14 = 21, overflow 1 
            ("0111", "1111", "0110", '1'),  -- 07 + 15 = 22, overflow 1 
            ("1000", "0000", "1000", '0'),  -- 08 + 00 = 08, overflow 0 
            ("1000", "0001", "1001", '0'),  -- 08 + 01 = 09, overflow 0 
            ("1000", "0010", "1010", '0'),  -- 08 + 02 = 10, overflow 0 
            ("1000", "0011", "1011", '0'),  -- 08 + 03 = 11, overflow 0 
            ("1000", "0100", "1100", '0'),  -- 08 + 04 = 12, overflow 0 
            ("1000", "0101", "1101", '0'),  -- 08 + 05 = 13, overflow 0 
            ("1000", "0110", "1110", '0'),  -- 08 + 06 = 14, overflow 0 
            ("1000", "0111", "1111", '0'),  -- 08 + 07 = 15, overflow 0 
            ("1000", "1000", "0000", '1'),  -- 08 + 08 = 16, overflow 1 
            ("1000", "1001", "0001", '1'),  -- 08 + 09 = 17, overflow 1 
            ("1000", "1010", "0010", '1'),  -- 08 + 10 = 18, overflow 1 
            ("1000", "1011", "0011", '1'),  -- 08 + 11 = 19, overflow 1 
            ("1000", "1100", "0100", '1'),  -- 08 + 12 = 20, overflow 1 
            ("1000", "1101", "0101", '1'),  -- 08 + 13 = 21, overflow 1 
            ("1000", "1110", "0110", '1'),  -- 08 + 14 = 22, overflow 1 
            ("1000", "1111", "0111", '1'),  -- 08 + 15 = 23, overflow 1 
            ("1001", "0000", "1001", '0'),  -- 09 + 00 = 09, overflow 0 
            ("1001", "0001", "1010", '0'),  -- 09 + 01 = 10, overflow 0 
            ("1001", "0010", "1011", '0'),  -- 09 + 02 = 11, overflow 0 
            ("1001", "0011", "1100", '0'),  -- 09 + 03 = 12, overflow 0 
            ("1001", "0100", "1101", '0'),  -- 09 + 04 = 13, overflow 0 
            ("1001", "0101", "1110", '0'),  -- 09 + 05 = 14, overflow 0 
            ("1001", "0110", "1111", '0'),  -- 09 + 06 = 15, overflow 0 
            ("1001", "0111", "0000", '1'),  -- 09 + 07 = 16, overflow 1 
            ("1001", "1000", "0001", '1'),  -- 09 + 08 = 17, overflow 1 
            ("1001", "1001", "0010", '1'),  -- 09 + 09 = 18, overflow 1 
            ("1001", "1010", "0011", '1'),  -- 09 + 10 = 19, overflow 1 
            ("1001", "1011", "0100", '1'),  -- 09 + 11 = 20, overflow 1 
            ("1001", "1100", "0101", '1'),  -- 09 + 12 = 21, overflow 1 
            ("1001", "1101", "0110", '1'),  -- 09 + 13 = 22, overflow 1 
            ("1001", "1110", "0111", '1'),  -- 09 + 14 = 23, overflow 1 
            ("1001", "1111", "1000", '1'),  -- 09 + 15 = 24, overflow 1 
            ("1010", "0000", "1010", '0'),  -- 10 + 00 = 10, overflow 0 
            ("1010", "0001", "1011", '0'),  -- 10 + 01 = 11, overflow 0 
            ("1010", "0010", "1100", '0'),  -- 10 + 02 = 12, overflow 0 
            ("1010", "0011", "1101", '0'),  -- 10 + 03 = 13, overflow 0 
            ("1010", "0100", "1110", '0'),  -- 10 + 04 = 14, overflow 0 
            ("1010", "0101", "1111", '0'),  -- 10 + 05 = 15, overflow 0 
            ("1010", "0110", "0000", '1'),  -- 10 + 06 = 16, overflow 1 
            ("1010", "0111", "0001", '1'),  -- 10 + 07 = 17, overflow 1 
            ("1010", "1000", "0010", '1'),  -- 10 + 08 = 18, overflow 1 
            ("1010", "1001", "0011", '1'),  -- 10 + 09 = 19, overflow 1 
            ("1010", "1010", "0100", '1'),  -- 10 + 10 = 20, overflow 1 
            ("1010", "1011", "0101", '1'),  -- 10 + 11 = 21, overflow 1 
            ("1010", "1100", "0110", '1'),  -- 10 + 12 = 22, overflow 1 
            ("1010", "1101", "0111", '1'),  -- 10 + 13 = 23, overflow 1 
            ("1010", "1110", "1000", '1'),  -- 10 + 14 = 24, overflow 1 
            ("1010", "1111", "1001", '1'),  -- 10 + 15 = 25, overflow 1 
            ("1011", "0000", "1011", '0'),  -- 11 + 00 = 11, overflow 0 
            ("1011", "0001", "1100", '0'),  -- 11 + 01 = 12, overflow 0 
            ("1011", "0010", "1101", '0'),  -- 11 + 02 = 13, overflow 0 
            ("1011", "0011", "1110", '0'),  -- 11 + 03 = 14, overflow 0 
            ("1011", "0100", "1111", '0'),  -- 11 + 04 = 15, overflow 0 
            ("1011", "0101", "0000", '1'),  -- 11 + 05 = 16, overflow 1 
            ("1011", "0110", "0001", '1'),  -- 11 + 06 = 17, overflow 1 
            ("1011", "0111", "0010", '1'),  -- 11 + 07 = 18, overflow 1 
            ("1011", "1000", "0011", '1'),  -- 11 + 08 = 19, overflow 1 
            ("1011", "1001", "0100", '1'),  -- 11 + 09 = 20, overflow 1 
            ("1011", "1010", "0101", '1'),  -- 11 + 10 = 21, overflow 1 
            ("1011", "1011", "0110", '1'),  -- 11 + 11 = 22, overflow 1 
            ("1011", "1100", "0111", '1'),  -- 11 + 12 = 23, overflow 1 
            ("1011", "1101", "1000", '1'),  -- 11 + 13 = 24, overflow 1 
            ("1011", "1110", "1001", '1'),  -- 11 + 14 = 25, overflow 1 
            ("1011", "1111", "1010", '1'),  -- 11 + 15 = 26, overflow 1 
            ("1100", "0000", "1100", '0'),  -- 12 + 00 = 12, overflow 0 
            ("1100", "0001", "1101", '0'),  -- 12 + 01 = 13, overflow 0 
            ("1100", "0010", "1110", '0'),  -- 12 + 02 = 14, overflow 0 
            ("1100", "0011", "1111", '0'),  -- 12 + 03 = 15, overflow 0 
            ("1100", "0100", "0000", '1'),  -- 12 + 04 = 16, overflow 1 
            ("1100", "0101", "0001", '1'),  -- 12 + 05 = 17, overflow 1 
            ("1100", "0110", "0010", '1'),  -- 12 + 06 = 18, overflow 1 
            ("1100", "0111", "0011", '1'),  -- 12 + 07 = 19, overflow 1 
            ("1100", "1000", "0100", '1'),  -- 12 + 08 = 20, overflow 1 
            ("1100", "1001", "0101", '1'),  -- 12 + 09 = 21, overflow 1 
            ("1100", "1010", "0110", '1'),  -- 12 + 10 = 22, overflow 1 
            ("1100", "1011", "0111", '1'),  -- 12 + 11 = 23, overflow 1 
            ("1100", "1100", "1000", '1'),  -- 12 + 12 = 24, overflow 1 
            ("1100", "1101", "1001", '1'),  -- 12 + 13 = 25, overflow 1 
            ("1100", "1110", "1010", '1'),  -- 12 + 14 = 26, overflow 1 
            ("1100", "1111", "1011", '1'),  -- 12 + 15 = 27, overflow 1 
            ("1101", "0000", "1101", '0'),  -- 13 + 00 = 13, overflow 0 
            ("1101", "0001", "1110", '0'),  -- 13 + 01 = 14, overflow 0 
            ("1101", "0010", "1111", '0'),  -- 13 + 02 = 15, overflow 0 
            ("1101", "0011", "0000", '1'),  -- 13 + 03 = 16, overflow 1 
            ("1101", "0100", "0001", '1'),  -- 13 + 04 = 17, overflow 1 
            ("1101", "0101", "0010", '1'),  -- 13 + 05 = 18, overflow 1 
            ("1101", "0110", "0011", '1'),  -- 13 + 06 = 19, overflow 1 
            ("1101", "0111", "0100", '1'),  -- 13 + 07 = 20, overflow 1 
            ("1101", "1000", "0101", '1'),  -- 13 + 08 = 21, overflow 1 
            ("1101", "1001", "0110", '1'),  -- 13 + 09 = 22, overflow 1 
            ("1101", "1010", "0111", '1'),  -- 13 + 10 = 23, overflow 1 
            ("1101", "1011", "1000", '1'),  -- 13 + 11 = 24, overflow 1 
            ("1101", "1100", "1001", '1'),  -- 13 + 12 = 25, overflow 1 
            ("1101", "1101", "1010", '1'),  -- 13 + 13 = 26, overflow 1 
            ("1101", "1110", "1011", '1'),  -- 13 + 14 = 27, overflow 1 
            ("1101", "1111", "1100", '1'),  -- 13 + 15 = 28, overflow 1 
            ("1110", "0000", "1110", '0'),  -- 14 + 00 = 14, overflow 0 
            ("1110", "0001", "1111", '0'),  -- 14 + 01 = 15, overflow 0 
            ("1110", "0010", "0000", '1'),  -- 14 + 02 = 16, overflow 1 
            ("1110", "0011", "0001", '1'),  -- 14 + 03 = 17, overflow 1 
            ("1110", "0100", "0010", '1'),  -- 14 + 04 = 18, overflow 1 
            ("1110", "0101", "0011", '1'),  -- 14 + 05 = 19, overflow 1 
            ("1110", "0110", "0100", '1'),  -- 14 + 06 = 20, overflow 1 
            ("1110", "0111", "0101", '1'),  -- 14 + 07 = 21, overflow 1 
            ("1110", "1000", "0110", '1'),  -- 14 + 08 = 22, overflow 1 
            ("1110", "1001", "0111", '1'),  -- 14 + 09 = 23, overflow 1 
            ("1110", "1010", "1000", '1'),  -- 14 + 10 = 24, overflow 1 
            ("1110", "1011", "1001", '1'),  -- 14 + 11 = 25, overflow 1 
            ("1110", "1100", "1010", '1'),  -- 14 + 12 = 26, overflow 1 
            ("1110", "1101", "1011", '1'),  -- 14 + 13 = 27, overflow 1 
            ("1110", "1110", "1100", '1'),  -- 14 + 14 = 28, overflow 1 
            ("1110", "1111", "1101", '1'),  -- 14 + 15 = 29, overflow 1 
            ("1111", "0000", "1111", '0'),  -- 15 + 00 = 15, overflow 0 
            ("1111", "0001", "0000", '1'),  -- 15 + 01 = 16, overflow 1 
            ("1111", "0010", "0001", '1'),  -- 15 + 02 = 17, overflow 1 
            ("1111", "0011", "0010", '1'),  -- 15 + 03 = 18, overflow 1 
            ("1111", "0100", "0011", '1'),  -- 15 + 04 = 19, overflow 1 
            ("1111", "0101", "0100", '1'),  -- 15 + 05 = 20, overflow 1 
            ("1111", "0110", "0101", '1'),  -- 15 + 06 = 21, overflow 1 
            ("1111", "0111", "0110", '1'),  -- 15 + 07 = 22, overflow 1 
            ("1111", "1000", "0111", '1'),  -- 15 + 08 = 23, overflow 1 
            ("1111", "1001", "1000", '1'),  -- 15 + 09 = 24, overflow 1 
            ("1111", "1010", "1001", '1'),  -- 15 + 10 = 25, overflow 1 
            ("1111", "1011", "1010", '1'),  -- 15 + 11 = 26, overflow 1 
            ("1111", "1100", "1011", '1'),  -- 15 + 12 = 27, overflow 1 
            ("1111", "1101", "1100", '1'),  -- 15 + 13 = 28, overflow 1 
            ("1111", "1110", "1101", '1'),  -- 15 + 14 = 29, overflow 1 
            ("1111", "1111", "1110", '1')   -- 15 + 15 = 30, overflow 1         
        );

    begin 

        for i in tabela_verdade'range loop
            
            -- entradas 
            a <= tabela_verdade(i).a;
            b <= tabela_verdade(i).b;

            -- espera os resultados
            wait for 1 ns;
            
            -- confere as saídas
            assert sum = tabela_verdade(i).sum report "Erro";
            assert cout = tabela_verdade(i).cout report "Erro";

        end loop;

        report "Fim dos teste";

        wait;

    end process;

end structural;